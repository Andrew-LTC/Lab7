`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/01/2021 09:16:18 PM
// Design Name: 
// Module Name: conseq_sequence
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module conseq_sequence(
    input clk,
    input reset_n,
    input x,
    output y
    );
    
    reg [2:0] state_reg, state_next;
    localparam s0 = 0;
    localparam s1 = 1;
    localparam s2 = 2;
    localparam s3 = 3;
    localparam s4 = 4;
    localparam s5 = 5;
    
    //State Register
    always @(posedge clk, negedge reset_n)
    begin
        if(~reset_n)
            state_reg <= s0;
        else
            state_reg <= state_next;
    end
    
    //Next State Logic
    always @(*)
    begin
        case(state_reg)
            s0: if(x)
                    state_next = s1;
                else
                    state_next = s2;
            s1: if(x)
                    state_next = s3;
                else
                    state_next = s0;
            s2: if(x)
                    state_next = s1;
                else
                    state_next = s4;
            s3: if(x)
                    state_next = s5;
                else
                    state_next = s0;
            s4: if(x)
                    state_next = s1;
                else
                    state_next = s4;
            s5: if(x)
                    state_next = s5;
                else
                    state_next = s0;
            default: state_next = state_reg;
        endcase
    end
    
    //Output Logic
    assign y = (state_reg == s4) | (state_reg == s5);
    
endmodule
